library verilog;
use verilog.vl_types.all;
entity cpu_vlg_tst is
end cpu_vlg_tst;
